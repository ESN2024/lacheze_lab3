library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
 
entity bcd_7segment is Port (
	bcd: in STD_LOGIC_VECTOR (3 downto 0);
	out7seg : out STD_LOGIC_VECTOR (7 downto 0));
end bcd_7segment;
 
architecture arch of bcd_7segment is
 
begin
 
 out7seg <= "11000000" when bcd = "0000" else
				"11111001" when bcd = "0001" else
            "10100100" when bcd = "0010" else
            "10110000" when bcd = "0011" else
            "10011001" when bcd = "0100" else
            "10010010" when bcd = "0101" else
            "10000010" when bcd = "0110" else
            "11111000" when bcd = "0111" else
            "10000000" when bcd = "1000" else
            "10010000" when bcd = "1001" else
				"10111111" when bcd = "1111" else
				"11111111";	
end architecture;
